-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"80cdac0c",
     3 => x"3a0b0b80",
     4 => x"c5ac0400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"80c5f32d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c4040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a7",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80cd",
   162 => x"98738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88aa0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0b8b",
   171 => x"a72d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0b8c",
   179 => x"d92d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80cda80c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"82c73f80",
   257 => x"c4ae3f04",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10101053",
   266 => x"51047381",
   267 => x"ff067383",
   268 => x"06098105",
   269 => x"83051010",
   270 => x"102b0772",
   271 => x"fc060c51",
   272 => x"51043c04",
   273 => x"72728072",
   274 => x"8106ff05",
   275 => x"09720605",
   276 => x"71105272",
   277 => x"0a100a53",
   278 => x"72ed3851",
   279 => x"51535104",
   280 => x"fe3d0d0b",
   281 => x"0b80dd94",
   282 => x"08538413",
   283 => x"0870882a",
   284 => x"70810651",
   285 => x"52527080",
   286 => x"2ef03871",
   287 => x"81ff0680",
   288 => x"0c843d0d",
   289 => x"04ff3d0d",
   290 => x"0b0b80dd",
   291 => x"94085271",
   292 => x"0870882a",
   293 => x"81327081",
   294 => x"06515151",
   295 => x"70f13873",
   296 => x"720c833d",
   297 => x"0d0480cd",
   298 => x"a808802e",
   299 => x"a43880cd",
   300 => x"ac08822e",
   301 => x"bd388380",
   302 => x"800b0b0b",
   303 => x"80dd940c",
   304 => x"82a0800b",
   305 => x"80dd980c",
   306 => x"8290800b",
   307 => x"80dd9c0c",
   308 => x"04f88080",
   309 => x"80a40b0b",
   310 => x"0b80dd94",
   311 => x"0cf88080",
   312 => x"82800b80",
   313 => x"dd980cf8",
   314 => x"80808480",
   315 => x"0b80dd9c",
   316 => x"0c0480c0",
   317 => x"a8808c0b",
   318 => x"0b0b80dd",
   319 => x"940c80c0",
   320 => x"a880940b",
   321 => x"80dd980c",
   322 => x"0b0b80cc",
   323 => x"e00b80dd",
   324 => x"9c0c04ff",
   325 => x"3d0d80dd",
   326 => x"a0335170",
   327 => x"a73880cd",
   328 => x"b4087008",
   329 => x"52527080",
   330 => x"2e943884",
   331 => x"1280cdb4",
   332 => x"0c702d80",
   333 => x"cdb40870",
   334 => x"08525270",
   335 => x"ee38810b",
   336 => x"80dda034",
   337 => x"833d0d04",
   338 => x"04803d0d",
   339 => x"0b0b80dd",
   340 => x"9008802e",
   341 => x"8e380b0b",
   342 => x"0b0b800b",
   343 => x"802e0981",
   344 => x"06853882",
   345 => x"3d0d040b",
   346 => x"0b80dd90",
   347 => x"510b0b0b",
   348 => x"f58e3f82",
   349 => x"3d0d0404",
   350 => x"fe3d0d89",
   351 => x"5380cce4",
   352 => x"5185f93f",
   353 => x"80ccf451",
   354 => x"85f23f81",
   355 => x"0a0b80dd",
   356 => x"ac0cff0b",
   357 => x"80ddb00c",
   358 => x"ff135372",
   359 => x"8025de38",
   360 => x"72800c84",
   361 => x"3d0d048c",
   362 => x"08028c0c",
   363 => x"f93d0d80",
   364 => x"0b8c08fc",
   365 => x"050c8c08",
   366 => x"88050880",
   367 => x"25ab388c",
   368 => x"08880508",
   369 => x"308c0888",
   370 => x"050c800b",
   371 => x"8c08f405",
   372 => x"0c8c08fc",
   373 => x"05088838",
   374 => x"810b8c08",
   375 => x"f4050c8c",
   376 => x"08f40508",
   377 => x"8c08fc05",
   378 => x"0c8c088c",
   379 => x"05088025",
   380 => x"ab388c08",
   381 => x"8c050830",
   382 => x"8c088c05",
   383 => x"0c800b8c",
   384 => x"08f0050c",
   385 => x"8c08fc05",
   386 => x"08883881",
   387 => x"0b8c08f0",
   388 => x"050c8c08",
   389 => x"f005088c",
   390 => x"08fc050c",
   391 => x"80538c08",
   392 => x"8c050852",
   393 => x"8c088805",
   394 => x"085181a7",
   395 => x"3f800870",
   396 => x"8c08f805",
   397 => x"0c548c08",
   398 => x"fc050880",
   399 => x"2e8c388c",
   400 => x"08f80508",
   401 => x"308c08f8",
   402 => x"050c8c08",
   403 => x"f8050870",
   404 => x"800c5489",
   405 => x"3d0d8c0c",
   406 => x"048c0802",
   407 => x"8c0cfb3d",
   408 => x"0d800b8c",
   409 => x"08fc050c",
   410 => x"8c088805",
   411 => x"08802593",
   412 => x"388c0888",
   413 => x"0508308c",
   414 => x"0888050c",
   415 => x"810b8c08",
   416 => x"fc050c8c",
   417 => x"088c0508",
   418 => x"80258c38",
   419 => x"8c088c05",
   420 => x"08308c08",
   421 => x"8c050c81",
   422 => x"538c088c",
   423 => x"0508528c",
   424 => x"08880508",
   425 => x"51ad3f80",
   426 => x"08708c08",
   427 => x"f8050c54",
   428 => x"8c08fc05",
   429 => x"08802e8c",
   430 => x"388c08f8",
   431 => x"0508308c",
   432 => x"08f8050c",
   433 => x"8c08f805",
   434 => x"0870800c",
   435 => x"54873d0d",
   436 => x"8c0c048c",
   437 => x"08028c0c",
   438 => x"fd3d0d81",
   439 => x"0b8c08fc",
   440 => x"050c800b",
   441 => x"8c08f805",
   442 => x"0c8c088c",
   443 => x"05088c08",
   444 => x"88050827",
   445 => x"ac388c08",
   446 => x"fc050880",
   447 => x"2ea33880",
   448 => x"0b8c088c",
   449 => x"05082499",
   450 => x"388c088c",
   451 => x"0508108c",
   452 => x"088c050c",
   453 => x"8c08fc05",
   454 => x"08108c08",
   455 => x"fc050cc9",
   456 => x"398c08fc",
   457 => x"0508802e",
   458 => x"80c9388c",
   459 => x"088c0508",
   460 => x"8c088805",
   461 => x"0826a138",
   462 => x"8c088805",
   463 => x"088c088c",
   464 => x"0508318c",
   465 => x"0888050c",
   466 => x"8c08f805",
   467 => x"088c08fc",
   468 => x"0508078c",
   469 => x"08f8050c",
   470 => x"8c08fc05",
   471 => x"08812a8c",
   472 => x"08fc050c",
   473 => x"8c088c05",
   474 => x"08812a8c",
   475 => x"088c050c",
   476 => x"ffaf398c",
   477 => x"08900508",
   478 => x"802e8f38",
   479 => x"8c088805",
   480 => x"08708c08",
   481 => x"f4050c51",
   482 => x"8d398c08",
   483 => x"f8050870",
   484 => x"8c08f405",
   485 => x"0c518c08",
   486 => x"f4050880",
   487 => x"0c853d0d",
   488 => x"8c0c04fc",
   489 => x"3d0d7670",
   490 => x"797b5555",
   491 => x"55558f72",
   492 => x"278c3872",
   493 => x"75078306",
   494 => x"5170802e",
   495 => x"a738ff12",
   496 => x"5271ff2e",
   497 => x"98387270",
   498 => x"81055433",
   499 => x"74708105",
   500 => x"5634ff12",
   501 => x"5271ff2e",
   502 => x"098106ea",
   503 => x"3874800c",
   504 => x"863d0d04",
   505 => x"74517270",
   506 => x"84055408",
   507 => x"71708405",
   508 => x"530c7270",
   509 => x"84055408",
   510 => x"71708405",
   511 => x"530c7270",
   512 => x"84055408",
   513 => x"71708405",
   514 => x"530c7270",
   515 => x"84055408",
   516 => x"71708405",
   517 => x"530cf012",
   518 => x"52718f26",
   519 => x"c9388372",
   520 => x"27953872",
   521 => x"70840554",
   522 => x"08717084",
   523 => x"05530cfc",
   524 => x"12527183",
   525 => x"26ed3870",
   526 => x"54ff8339",
   527 => x"f73d0d7c",
   528 => x"70525380",
   529 => x"c83f7254",
   530 => x"80085580",
   531 => x"cd845681",
   532 => x"57800881",
   533 => x"055a8b3d",
   534 => x"e4115953",
   535 => x"8259f413",
   536 => x"527b8811",
   537 => x"08525381",
   538 => x"833f8008",
   539 => x"30708008",
   540 => x"079f2c8a",
   541 => x"07800c53",
   542 => x"8b3d0d04",
   543 => x"ff3d0d73",
   544 => x"5280cdb8",
   545 => x"0851ffb4",
   546 => x"3f833d0d",
   547 => x"04fd3d0d",
   548 => x"75707183",
   549 => x"06535552",
   550 => x"70b83871",
   551 => x"70087009",
   552 => x"f7fbfdff",
   553 => x"120670f8",
   554 => x"84828180",
   555 => x"06515152",
   556 => x"53709d38",
   557 => x"84137008",
   558 => x"7009f7fb",
   559 => x"fdff1206",
   560 => x"70f88482",
   561 => x"81800651",
   562 => x"51525370",
   563 => x"802ee538",
   564 => x"72527133",
   565 => x"5170802e",
   566 => x"8a388112",
   567 => x"70335252",
   568 => x"70f83871",
   569 => x"7431800c",
   570 => x"853d0d04",
   571 => x"f23d0d60",
   572 => x"62881108",
   573 => x"7057575f",
   574 => x"5a74802e",
   575 => x"8190388c",
   576 => x"1a227083",
   577 => x"2a813270",
   578 => x"81065155",
   579 => x"58738638",
   580 => x"901a0891",
   581 => x"38795190",
   582 => x"a23fff54",
   583 => x"800880ee",
   584 => x"388c1a22",
   585 => x"587d0857",
   586 => x"807883ff",
   587 => x"ff06700a",
   588 => x"100a7081",
   589 => x"06515657",
   590 => x"5573752e",
   591 => x"80d73874",
   592 => x"90387608",
   593 => x"84180888",
   594 => x"19595659",
   595 => x"74802ef2",
   596 => x"38745488",
   597 => x"80752784",
   598 => x"38888054",
   599 => x"73537852",
   600 => x"9c1a0851",
   601 => x"a41a0854",
   602 => x"732d800b",
   603 => x"80082582",
   604 => x"e6388008",
   605 => x"19758008",
   606 => x"317f8805",
   607 => x"08800831",
   608 => x"70618805",
   609 => x"0c565659",
   610 => x"73ffb438",
   611 => x"80547380",
   612 => x"0c903d0d",
   613 => x"04758132",
   614 => x"70810676",
   615 => x"41515473",
   616 => x"802e81c1",
   617 => x"38749038",
   618 => x"76088418",
   619 => x"08881959",
   620 => x"56597480",
   621 => x"2ef23888",
   622 => x"1a087883",
   623 => x"ffff0670",
   624 => x"892a7081",
   625 => x"06515659",
   626 => x"5673802e",
   627 => x"82fa3875",
   628 => x"75278d38",
   629 => x"77872a70",
   630 => x"81065154",
   631 => x"7382b538",
   632 => x"74762783",
   633 => x"38745675",
   634 => x"53785279",
   635 => x"08518582",
   636 => x"3f881a08",
   637 => x"7631881b",
   638 => x"0c790816",
   639 => x"7a0c7456",
   640 => x"75197577",
   641 => x"317f8805",
   642 => x"08783170",
   643 => x"6188050c",
   644 => x"56565973",
   645 => x"802efef4",
   646 => x"388c1a22",
   647 => x"58ff8639",
   648 => x"77785479",
   649 => x"537b5256",
   650 => x"84c83f88",
   651 => x"1a087831",
   652 => x"881b0c79",
   653 => x"08187a0c",
   654 => x"7c76315d",
   655 => x"7c8e3879",
   656 => x"518fdc3f",
   657 => x"8008818f",
   658 => x"3880085f",
   659 => x"75197577",
   660 => x"317f8805",
   661 => x"08783170",
   662 => x"6188050c",
   663 => x"56565973",
   664 => x"802efea8",
   665 => x"38748183",
   666 => x"38760884",
   667 => x"18088819",
   668 => x"59565974",
   669 => x"802ef238",
   670 => x"74538a52",
   671 => x"785182d3",
   672 => x"3f800879",
   673 => x"3181055d",
   674 => x"80088438",
   675 => x"81155d81",
   676 => x"5f7c5874",
   677 => x"7d278338",
   678 => x"7458941a",
   679 => x"08881b08",
   680 => x"11575c80",
   681 => x"7a085c54",
   682 => x"901a087b",
   683 => x"27833881",
   684 => x"54757825",
   685 => x"843873ba",
   686 => x"387b7824",
   687 => x"fee2387b",
   688 => x"5378529c",
   689 => x"1a0851a4",
   690 => x"1a085473",
   691 => x"2d800856",
   692 => x"80088024",
   693 => x"fee2388c",
   694 => x"1a2280c0",
   695 => x"0754738c",
   696 => x"1b23ff54",
   697 => x"73800c90",
   698 => x"3d0d047e",
   699 => x"ffa338ff",
   700 => x"87397553",
   701 => x"78527a51",
   702 => x"82f83f79",
   703 => x"08167a0c",
   704 => x"79518e9b",
   705 => x"3f8008cf",
   706 => x"387c7631",
   707 => x"5d7cfebc",
   708 => x"38feac39",
   709 => x"901a087a",
   710 => x"08713176",
   711 => x"1170565a",
   712 => x"575280cd",
   713 => x"b8085184",
   714 => x"8c3f8008",
   715 => x"802effa7",
   716 => x"38800890",
   717 => x"1b0c8008",
   718 => x"167a0c77",
   719 => x"941b0c74",
   720 => x"881b0c74",
   721 => x"56fd9939",
   722 => x"79085890",
   723 => x"1a087827",
   724 => x"83388154",
   725 => x"75752784",
   726 => x"3873b338",
   727 => x"941a0856",
   728 => x"75752680",
   729 => x"d3387553",
   730 => x"78529c1a",
   731 => x"0851a41a",
   732 => x"0854732d",
   733 => x"80085680",
   734 => x"088024fd",
   735 => x"83388c1a",
   736 => x"2280c007",
   737 => x"54738c1b",
   738 => x"23ff54fe",
   739 => x"d7397553",
   740 => x"78527751",
   741 => x"81dc3f79",
   742 => x"08167a0c",
   743 => x"79518cff",
   744 => x"3f800880",
   745 => x"2efcd938",
   746 => x"8c1a2280",
   747 => x"c0075473",
   748 => x"8c1b23ff",
   749 => x"54fead39",
   750 => x"74755479",
   751 => x"53785256",
   752 => x"81b03f88",
   753 => x"1a087531",
   754 => x"881b0c79",
   755 => x"08157a0c",
   756 => x"fcae39fa",
   757 => x"3d0d7a79",
   758 => x"028805a7",
   759 => x"05335652",
   760 => x"53837327",
   761 => x"8a387083",
   762 => x"06527180",
   763 => x"2ea838ff",
   764 => x"135372ff",
   765 => x"2e973870",
   766 => x"33527372",
   767 => x"2e913881",
   768 => x"11ff1454",
   769 => x"5172ff2e",
   770 => x"098106eb",
   771 => x"38805170",
   772 => x"800c883d",
   773 => x"0d047072",
   774 => x"57558351",
   775 => x"75828029",
   776 => x"14ff1252",
   777 => x"56708025",
   778 => x"f3388373",
   779 => x"27bf3874",
   780 => x"08763270",
   781 => x"09f7fbfd",
   782 => x"ff120670",
   783 => x"f8848281",
   784 => x"80065151",
   785 => x"5170802e",
   786 => x"99387451",
   787 => x"80527033",
   788 => x"5773772e",
   789 => x"ffb93881",
   790 => x"11811353",
   791 => x"51837227",
   792 => x"ed38fc13",
   793 => x"84165653",
   794 => x"728326c3",
   795 => x"387451fe",
   796 => x"fe39fa3d",
   797 => x"0d787a7c",
   798 => x"72727257",
   799 => x"57575956",
   800 => x"56747627",
   801 => x"b2387615",
   802 => x"51757127",
   803 => x"aa387077",
   804 => x"17ff1454",
   805 => x"555371ff",
   806 => x"2e9638ff",
   807 => x"14ff1454",
   808 => x"54723374",
   809 => x"34ff1252",
   810 => x"71ff2e09",
   811 => x"8106ec38",
   812 => x"75800c88",
   813 => x"3d0d0476",
   814 => x"8f269738",
   815 => x"ff125271",
   816 => x"ff2eed38",
   817 => x"72708105",
   818 => x"54337470",
   819 => x"81055634",
   820 => x"eb397476",
   821 => x"07830651",
   822 => x"70e23875",
   823 => x"75545172",
   824 => x"70840554",
   825 => x"08717084",
   826 => x"05530c72",
   827 => x"70840554",
   828 => x"08717084",
   829 => x"05530c72",
   830 => x"70840554",
   831 => x"08717084",
   832 => x"05530c72",
   833 => x"70840554",
   834 => x"08717084",
   835 => x"05530cf0",
   836 => x"1252718f",
   837 => x"26c93883",
   838 => x"72279538",
   839 => x"72708405",
   840 => x"54087170",
   841 => x"8405530c",
   842 => x"fc125271",
   843 => x"8326ed38",
   844 => x"7054ff88",
   845 => x"39ef3d0d",
   846 => x"63656740",
   847 => x"5d427b80",
   848 => x"2e84fa38",
   849 => x"6151a5b6",
   850 => x"3ff81c70",
   851 => x"84120870",
   852 => x"fc067062",
   853 => x"8b0570f8",
   854 => x"06415945",
   855 => x"5b5c4157",
   856 => x"96742782",
   857 => x"c338807b",
   858 => x"247e7c26",
   859 => x"07598054",
   860 => x"78742e09",
   861 => x"810682a9",
   862 => x"38777b25",
   863 => x"81fc3877",
   864 => x"1780d4f4",
   865 => x"0b880508",
   866 => x"5e567c76",
   867 => x"2e84bd38",
   868 => x"84160870",
   869 => x"fe061784",
   870 => x"11088106",
   871 => x"51555573",
   872 => x"828b3874",
   873 => x"fc06597c",
   874 => x"762e84dd",
   875 => x"3877195f",
   876 => x"7e7b2581",
   877 => x"fd387981",
   878 => x"06547382",
   879 => x"bf387677",
   880 => x"08318411",
   881 => x"08fc0656",
   882 => x"5a75802e",
   883 => x"91387c76",
   884 => x"2e84ea38",
   885 => x"74191859",
   886 => x"787b2584",
   887 => x"89387980",
   888 => x"2e829938",
   889 => x"7715567a",
   890 => x"76248290",
   891 => x"388c1a08",
   892 => x"881b0871",
   893 => x"8c120c88",
   894 => x"120c5579",
   895 => x"76595788",
   896 => x"1761fc05",
   897 => x"575975a4",
   898 => x"2685ef38",
   899 => x"7b795555",
   900 => x"93762780",
   901 => x"c9387b70",
   902 => x"84055d08",
   903 => x"7c56790c",
   904 => x"74708405",
   905 => x"56088c18",
   906 => x"0c901754",
   907 => x"9b7627ae",
   908 => x"38747084",
   909 => x"05560874",
   910 => x"0c747084",
   911 => x"05560894",
   912 => x"180c9817",
   913 => x"54a37627",
   914 => x"95387470",
   915 => x"84055608",
   916 => x"740c7470",
   917 => x"84055608",
   918 => x"9c180ca0",
   919 => x"17547470",
   920 => x"84055608",
   921 => x"74708405",
   922 => x"560c7470",
   923 => x"84055608",
   924 => x"74708405",
   925 => x"560c7408",
   926 => x"740c777b",
   927 => x"3156758f",
   928 => x"2680c938",
   929 => x"84170881",
   930 => x"06780784",
   931 => x"180c7717",
   932 => x"84110881",
   933 => x"0784120c",
   934 => x"546151a2",
   935 => x"e23f8817",
   936 => x"5473800c",
   937 => x"933d0d04",
   938 => x"905bfdba",
   939 => x"397856fe",
   940 => x"85398c16",
   941 => x"08881708",
   942 => x"718c120c",
   943 => x"88120c55",
   944 => x"7e707c31",
   945 => x"57588f76",
   946 => x"27ffb938",
   947 => x"7a178418",
   948 => x"0881067c",
   949 => x"0784190c",
   950 => x"76810784",
   951 => x"120c7611",
   952 => x"84110881",
   953 => x"0784120c",
   954 => x"55880552",
   955 => x"61518cf7",
   956 => x"3f6151a2",
   957 => x"8a3f8817",
   958 => x"54ffa639",
   959 => x"7d526151",
   960 => x"94f73f80",
   961 => x"08598008",
   962 => x"802e81a3",
   963 => x"388008f8",
   964 => x"05608405",
   965 => x"08fe0661",
   966 => x"05555776",
   967 => x"742e83e6",
   968 => x"38fc1856",
   969 => x"75a42681",
   970 => x"aa387b80",
   971 => x"08555593",
   972 => x"762780d8",
   973 => x"38747084",
   974 => x"05560880",
   975 => x"08708405",
   976 => x"800c0c80",
   977 => x"08757084",
   978 => x"05570871",
   979 => x"70840553",
   980 => x"0c549b76",
   981 => x"27b63874",
   982 => x"70840556",
   983 => x"08747084",
   984 => x"05560c74",
   985 => x"70840556",
   986 => x"08747084",
   987 => x"05560ca3",
   988 => x"76279938",
   989 => x"74708405",
   990 => x"56087470",
   991 => x"8405560c",
   992 => x"74708405",
   993 => x"56087470",
   994 => x"8405560c",
   995 => x"74708405",
   996 => x"56087470",
   997 => x"8405560c",
   998 => x"74708405",
   999 => x"56087470",
  1000 => x"8405560c",
  1001 => x"7408740c",
  1002 => x"7b526151",
  1003 => x"8bb93f61",
  1004 => x"51a0cc3f",
  1005 => x"78547380",
  1006 => x"0c933d0d",
  1007 => x"047d5261",
  1008 => x"5193b63f",
  1009 => x"8008800c",
  1010 => x"933d0d04",
  1011 => x"84160855",
  1012 => x"fbd13975",
  1013 => x"537b5280",
  1014 => x"0851efc7",
  1015 => x"3f7b5261",
  1016 => x"518b843f",
  1017 => x"ca398c16",
  1018 => x"08881708",
  1019 => x"718c120c",
  1020 => x"88120c55",
  1021 => x"8c1a0888",
  1022 => x"1b08718c",
  1023 => x"120c8812",
  1024 => x"0c557979",
  1025 => x"5957fbf7",
  1026 => x"39771990",
  1027 => x"1c555573",
  1028 => x"7524fba2",
  1029 => x"387a1770",
  1030 => x"80d4f40b",
  1031 => x"88050c75",
  1032 => x"7c318107",
  1033 => x"84120c5d",
  1034 => x"84170881",
  1035 => x"067b0784",
  1036 => x"180c6151",
  1037 => x"9fc93f88",
  1038 => x"1754fce5",
  1039 => x"39741918",
  1040 => x"901c555d",
  1041 => x"737d24fb",
  1042 => x"95388c1a",
  1043 => x"08881b08",
  1044 => x"718c120c",
  1045 => x"88120c55",
  1046 => x"881a61fc",
  1047 => x"05575975",
  1048 => x"a42681ae",
  1049 => x"387b7955",
  1050 => x"55937627",
  1051 => x"80c9387b",
  1052 => x"7084055d",
  1053 => x"087c5679",
  1054 => x"0c747084",
  1055 => x"0556088c",
  1056 => x"1b0c901a",
  1057 => x"549b7627",
  1058 => x"ae387470",
  1059 => x"84055608",
  1060 => x"740c7470",
  1061 => x"84055608",
  1062 => x"941b0c98",
  1063 => x"1a54a376",
  1064 => x"27953874",
  1065 => x"70840556",
  1066 => x"08740c74",
  1067 => x"70840556",
  1068 => x"089c1b0c",
  1069 => x"a01a5474",
  1070 => x"70840556",
  1071 => x"08747084",
  1072 => x"05560c74",
  1073 => x"70840556",
  1074 => x"08747084",
  1075 => x"05560c74",
  1076 => x"08740c7a",
  1077 => x"1a7080d4",
  1078 => x"f40b8805",
  1079 => x"0c7d7c31",
  1080 => x"81078412",
  1081 => x"0c54841a",
  1082 => x"0881067b",
  1083 => x"07841b0c",
  1084 => x"61519e8b",
  1085 => x"3f7854fd",
  1086 => x"bd397553",
  1087 => x"7b527851",
  1088 => x"eda13ffa",
  1089 => x"f5398417",
  1090 => x"08fc0618",
  1091 => x"605858fa",
  1092 => x"e9397553",
  1093 => x"7b527851",
  1094 => x"ed893f7a",
  1095 => x"1a7080d4",
  1096 => x"f40b8805",
  1097 => x"0c7d7c31",
  1098 => x"81078412",
  1099 => x"0c54841a",
  1100 => x"0881067b",
  1101 => x"07841b0c",
  1102 => x"ffb639fa",
  1103 => x"3d0d7880",
  1104 => x"cdb80854",
  1105 => x"55b81308",
  1106 => x"802e81b6",
  1107 => x"388c1522",
  1108 => x"7083ffff",
  1109 => x"0670832a",
  1110 => x"81327081",
  1111 => x"06515555",
  1112 => x"5672802e",
  1113 => x"80dc3873",
  1114 => x"842a8132",
  1115 => x"810657ff",
  1116 => x"537680f7",
  1117 => x"3873822a",
  1118 => x"70810651",
  1119 => x"5372802e",
  1120 => x"b938b015",
  1121 => x"08547380",
  1122 => x"2e9c3880",
  1123 => x"c0155373",
  1124 => x"732e8f38",
  1125 => x"735280cd",
  1126 => x"b8085187",
  1127 => x"ca3f8c15",
  1128 => x"225676b0",
  1129 => x"160c75db",
  1130 => x"0653728c",
  1131 => x"1623800b",
  1132 => x"84160c90",
  1133 => x"1508750c",
  1134 => x"72567588",
  1135 => x"0753728c",
  1136 => x"16239015",
  1137 => x"08802e80",
  1138 => x"c1388c15",
  1139 => x"22708106",
  1140 => x"5553739e",
  1141 => x"38720a10",
  1142 => x"0a708106",
  1143 => x"51537285",
  1144 => x"38941508",
  1145 => x"54738816",
  1146 => x"0c805372",
  1147 => x"800c883d",
  1148 => x"0d04800b",
  1149 => x"88160c94",
  1150 => x"15083098",
  1151 => x"160c8053",
  1152 => x"ea397251",
  1153 => x"82fb3ffe",
  1154 => x"c4397451",
  1155 => x"8ce83f8c",
  1156 => x"15227081",
  1157 => x"06555373",
  1158 => x"802effb9",
  1159 => x"38d439f8",
  1160 => x"3d0d7a58",
  1161 => x"77802e81",
  1162 => x"993880cd",
  1163 => x"b80854b8",
  1164 => x"1408802e",
  1165 => x"80ed388c",
  1166 => x"18227090",
  1167 => x"2b70902c",
  1168 => x"70832a81",
  1169 => x"3281065c",
  1170 => x"51575478",
  1171 => x"80cd3890",
  1172 => x"18085776",
  1173 => x"802e80c3",
  1174 => x"38770877",
  1175 => x"3177790c",
  1176 => x"7683067a",
  1177 => x"58555573",
  1178 => x"85389418",
  1179 => x"08567588",
  1180 => x"190c8075",
  1181 => x"25a53874",
  1182 => x"5376529c",
  1183 => x"180851a4",
  1184 => x"18085473",
  1185 => x"2d800b80",
  1186 => x"082580c9",
  1187 => x"38800817",
  1188 => x"75800831",
  1189 => x"56577480",
  1190 => x"24dd3880",
  1191 => x"0b800c8a",
  1192 => x"3d0d0473",
  1193 => x"5181da3f",
  1194 => x"8c182270",
  1195 => x"902b7090",
  1196 => x"2c70832a",
  1197 => x"81328106",
  1198 => x"5c515754",
  1199 => x"78dd38ff",
  1200 => x"8e39a49f",
  1201 => x"5280cdb8",
  1202 => x"085189f1",
  1203 => x"3f800880",
  1204 => x"0c8a3d0d",
  1205 => x"048c1822",
  1206 => x"80c00754",
  1207 => x"738c1923",
  1208 => x"ff0b800c",
  1209 => x"8a3d0d04",
  1210 => x"803d0d72",
  1211 => x"5180710c",
  1212 => x"800b8412",
  1213 => x"0c800b88",
  1214 => x"120c028e",
  1215 => x"05228c12",
  1216 => x"23029205",
  1217 => x"228e1223",
  1218 => x"800b9012",
  1219 => x"0c800b94",
  1220 => x"120c800b",
  1221 => x"98120c70",
  1222 => x"9c120c80",
  1223 => x"c0b40ba0",
  1224 => x"120c80c1",
  1225 => x"800ba412",
  1226 => x"0c80c1fc",
  1227 => x"0ba8120c",
  1228 => x"80c2cd0b",
  1229 => x"ac120c82",
  1230 => x"3d0d04fa",
  1231 => x"3d0d7970",
  1232 => x"80dc298c",
  1233 => x"11547a53",
  1234 => x"56578cad",
  1235 => x"3f800880",
  1236 => x"08555680",
  1237 => x"08802ea2",
  1238 => x"3880088c",
  1239 => x"0554800b",
  1240 => x"80080c76",
  1241 => x"80088405",
  1242 => x"0c738008",
  1243 => x"88050c74",
  1244 => x"53805273",
  1245 => x"5197f83f",
  1246 => x"75547380",
  1247 => x"0c883d0d",
  1248 => x"04fc3d0d",
  1249 => x"76a9940b",
  1250 => x"bc120c55",
  1251 => x"810bb816",
  1252 => x"0c800b84",
  1253 => x"dc160c83",
  1254 => x"0b84e016",
  1255 => x"0c84e815",
  1256 => x"84e4160c",
  1257 => x"74548053",
  1258 => x"84528415",
  1259 => x"0851feb8",
  1260 => x"3f745481",
  1261 => x"53895288",
  1262 => x"150851fe",
  1263 => x"ab3f7454",
  1264 => x"82538a52",
  1265 => x"8c150851",
  1266 => x"fe9e3f86",
  1267 => x"3d0d04f9",
  1268 => x"3d0d7980",
  1269 => x"cdb80854",
  1270 => x"57b81308",
  1271 => x"802e80c8",
  1272 => x"3884dc13",
  1273 => x"56881608",
  1274 => x"841708ff",
  1275 => x"05555580",
  1276 => x"74249f38",
  1277 => x"8c152270",
  1278 => x"902b7090",
  1279 => x"2c515458",
  1280 => x"72802e80",
  1281 => x"ca3880dc",
  1282 => x"15ff1555",
  1283 => x"55738025",
  1284 => x"e3387508",
  1285 => x"5372802e",
  1286 => x"9f387256",
  1287 => x"88160884",
  1288 => x"1708ff05",
  1289 => x"5555c839",
  1290 => x"7251fed5",
  1291 => x"3f80cdb8",
  1292 => x"0884dc05",
  1293 => x"56ffae39",
  1294 => x"84527651",
  1295 => x"fdfd3f80",
  1296 => x"08760c80",
  1297 => x"08802e80",
  1298 => x"c0388008",
  1299 => x"56ce3981",
  1300 => x"0b8c1623",
  1301 => x"72750c72",
  1302 => x"88160c72",
  1303 => x"84160c72",
  1304 => x"90160c72",
  1305 => x"94160c72",
  1306 => x"98160cff",
  1307 => x"0b8e1623",
  1308 => x"72b0160c",
  1309 => x"72b4160c",
  1310 => x"7280c416",
  1311 => x"0c7280c8",
  1312 => x"160c7480",
  1313 => x"0c893d0d",
  1314 => x"048c770c",
  1315 => x"800b800c",
  1316 => x"893d0d04",
  1317 => x"ff3d0da4",
  1318 => x"9f527351",
  1319 => x"869f3f83",
  1320 => x"3d0d0480",
  1321 => x"3d0d80cd",
  1322 => x"b80851e8",
  1323 => x"3f823d0d",
  1324 => x"04fb3d0d",
  1325 => x"77705256",
  1326 => x"96c43f80",
  1327 => x"d4f40b88",
  1328 => x"05088411",
  1329 => x"08fc0670",
  1330 => x"7b319fef",
  1331 => x"05e08006",
  1332 => x"e0800556",
  1333 => x"5653a080",
  1334 => x"74249438",
  1335 => x"80527551",
  1336 => x"969e3f80",
  1337 => x"d4fc0815",
  1338 => x"53728008",
  1339 => x"2e8f3875",
  1340 => x"51968c3f",
  1341 => x"80537280",
  1342 => x"0c873d0d",
  1343 => x"04733052",
  1344 => x"755195fc",
  1345 => x"3f8008ff",
  1346 => x"2ea83880",
  1347 => x"d4f40b88",
  1348 => x"05087575",
  1349 => x"31810784",
  1350 => x"120c5380",
  1351 => x"d4b80874",
  1352 => x"3180d4b8",
  1353 => x"0c755195",
  1354 => x"d63f810b",
  1355 => x"800c873d",
  1356 => x"0d048052",
  1357 => x"755195c8",
  1358 => x"3f80d4f4",
  1359 => x"0b880508",
  1360 => x"80087131",
  1361 => x"56538f75",
  1362 => x"25ffa438",
  1363 => x"800880d4",
  1364 => x"e8083180",
  1365 => x"d4b80c74",
  1366 => x"81078414",
  1367 => x"0c755195",
  1368 => x"9e3f8053",
  1369 => x"ff9039f6",
  1370 => x"3d0d7c7e",
  1371 => x"545b7280",
  1372 => x"2e828338",
  1373 => x"7a519586",
  1374 => x"3ff81384",
  1375 => x"110870fe",
  1376 => x"06701384",
  1377 => x"1108fc06",
  1378 => x"5d585954",
  1379 => x"5880d4fc",
  1380 => x"08752e82",
  1381 => x"de387884",
  1382 => x"160c8073",
  1383 => x"8106545a",
  1384 => x"727a2e81",
  1385 => x"d5387815",
  1386 => x"84110881",
  1387 => x"06515372",
  1388 => x"a0387817",
  1389 => x"577981e6",
  1390 => x"38881508",
  1391 => x"537280d4",
  1392 => x"fc2e82f9",
  1393 => x"388c1508",
  1394 => x"708c150c",
  1395 => x"7388120c",
  1396 => x"56768107",
  1397 => x"84190c76",
  1398 => x"1877710c",
  1399 => x"53798191",
  1400 => x"3883ff77",
  1401 => x"2781c838",
  1402 => x"76892a77",
  1403 => x"832a5653",
  1404 => x"72802ebf",
  1405 => x"3876862a",
  1406 => x"b8055584",
  1407 => x"7327b438",
  1408 => x"80db1355",
  1409 => x"947327ab",
  1410 => x"38768c2a",
  1411 => x"80ee0555",
  1412 => x"80d47327",
  1413 => x"9e38768f",
  1414 => x"2a80f705",
  1415 => x"5582d473",
  1416 => x"27913876",
  1417 => x"922a80fc",
  1418 => x"05558ad4",
  1419 => x"73278438",
  1420 => x"80fe5574",
  1421 => x"10101080",
  1422 => x"d4f40588",
  1423 => x"11085556",
  1424 => x"73762e82",
  1425 => x"b3388414",
  1426 => x"08fc0653",
  1427 => x"7673278d",
  1428 => x"38881408",
  1429 => x"5473762e",
  1430 => x"098106ea",
  1431 => x"388c1408",
  1432 => x"708c1a0c",
  1433 => x"74881a0c",
  1434 => x"7888120c",
  1435 => x"56778c15",
  1436 => x"0c7a5193",
  1437 => x"8a3f8c3d",
  1438 => x"0d047708",
  1439 => x"78713159",
  1440 => x"77058819",
  1441 => x"08545772",
  1442 => x"80d4fc2e",
  1443 => x"80e0388c",
  1444 => x"1808708c",
  1445 => x"150c7388",
  1446 => x"120c56fe",
  1447 => x"89398815",
  1448 => x"088c1608",
  1449 => x"708c130c",
  1450 => x"5788170c",
  1451 => x"fea33976",
  1452 => x"832a7054",
  1453 => x"55807524",
  1454 => x"81983872",
  1455 => x"822c8171",
  1456 => x"2b80d4f8",
  1457 => x"080780d4",
  1458 => x"f40b8405",
  1459 => x"0c537410",
  1460 => x"101080d4",
  1461 => x"f4058811",
  1462 => x"08555675",
  1463 => x"8c190c73",
  1464 => x"88190c77",
  1465 => x"88170c77",
  1466 => x"8c150cff",
  1467 => x"8439815a",
  1468 => x"fdb43978",
  1469 => x"17738106",
  1470 => x"54577298",
  1471 => x"38770878",
  1472 => x"71315977",
  1473 => x"058c1908",
  1474 => x"881a0871",
  1475 => x"8c120c88",
  1476 => x"120c5757",
  1477 => x"76810784",
  1478 => x"190c7780",
  1479 => x"d4f40b88",
  1480 => x"050c80d4",
  1481 => x"f0087726",
  1482 => x"fec73880",
  1483 => x"d4ec0852",
  1484 => x"7a51fafd",
  1485 => x"3f7a5191",
  1486 => x"c63ffeba",
  1487 => x"3981788c",
  1488 => x"150c7888",
  1489 => x"150c738c",
  1490 => x"1a0c7388",
  1491 => x"1a0c5afd",
  1492 => x"80398315",
  1493 => x"70822c81",
  1494 => x"712b80d4",
  1495 => x"f8080780",
  1496 => x"d4f40b84",
  1497 => x"050c5153",
  1498 => x"74101010",
  1499 => x"80d4f405",
  1500 => x"88110855",
  1501 => x"56fee439",
  1502 => x"74538075",
  1503 => x"24a73872",
  1504 => x"822c8171",
  1505 => x"2b80d4f8",
  1506 => x"080780d4",
  1507 => x"f40b8405",
  1508 => x"0c53758c",
  1509 => x"190c7388",
  1510 => x"190c7788",
  1511 => x"170c778c",
  1512 => x"150cfdcd",
  1513 => x"39831570",
  1514 => x"822c8171",
  1515 => x"2b80d4f8",
  1516 => x"080780d4",
  1517 => x"f40b8405",
  1518 => x"0c5153d6",
  1519 => x"39f93d0d",
  1520 => x"797b5853",
  1521 => x"800b80cd",
  1522 => x"b8085356",
  1523 => x"72722e80",
  1524 => x"c03884dc",
  1525 => x"13557476",
  1526 => x"2eb73888",
  1527 => x"15088416",
  1528 => x"08ff0554",
  1529 => x"54807324",
  1530 => x"9d388c14",
  1531 => x"2270902b",
  1532 => x"70902c51",
  1533 => x"53587180",
  1534 => x"d83880dc",
  1535 => x"14ff1454",
  1536 => x"54728025",
  1537 => x"e5387408",
  1538 => x"5574d038",
  1539 => x"80cdb808",
  1540 => x"5284dc12",
  1541 => x"5574802e",
  1542 => x"b1388815",
  1543 => x"08841608",
  1544 => x"ff055454",
  1545 => x"8073249c",
  1546 => x"388c1422",
  1547 => x"70902b70",
  1548 => x"902c5153",
  1549 => x"5871ad38",
  1550 => x"80dc14ff",
  1551 => x"14545472",
  1552 => x"8025e638",
  1553 => x"74085574",
  1554 => x"d1387580",
  1555 => x"0c893d0d",
  1556 => x"04735176",
  1557 => x"2d758008",
  1558 => x"0780dc15",
  1559 => x"ff155555",
  1560 => x"56ff9e39",
  1561 => x"7351762d",
  1562 => x"75800807",
  1563 => x"80dc15ff",
  1564 => x"15555556",
  1565 => x"ca39ea3d",
  1566 => x"0d688c11",
  1567 => x"22700a10",
  1568 => x"0a810657",
  1569 => x"58567480",
  1570 => x"e4388e16",
  1571 => x"2270902b",
  1572 => x"70902c51",
  1573 => x"55588074",
  1574 => x"24b13898",
  1575 => x"3dc40553",
  1576 => x"735280cd",
  1577 => x"b8085192",
  1578 => x"ac3f800b",
  1579 => x"80082497",
  1580 => x"387983e0",
  1581 => x"80065473",
  1582 => x"80c0802e",
  1583 => x"818f3873",
  1584 => x"8280802e",
  1585 => x"8191388c",
  1586 => x"16225776",
  1587 => x"90800754",
  1588 => x"738c1723",
  1589 => x"88805280",
  1590 => x"cdb80851",
  1591 => x"819b3f80",
  1592 => x"089d388c",
  1593 => x"16228207",
  1594 => x"54738c17",
  1595 => x"2380c316",
  1596 => x"70770c90",
  1597 => x"170c810b",
  1598 => x"94170c98",
  1599 => x"3d0d0480",
  1600 => x"cdb808a9",
  1601 => x"940bbc12",
  1602 => x"0c548c16",
  1603 => x"22818007",
  1604 => x"54738c17",
  1605 => x"23800876",
  1606 => x"0c800890",
  1607 => x"170c8880",
  1608 => x"0b94170c",
  1609 => x"74802ed3",
  1610 => x"388e1622",
  1611 => x"70902b70",
  1612 => x"902c5355",
  1613 => x"5898a23f",
  1614 => x"8008802e",
  1615 => x"ffbd388c",
  1616 => x"16228107",
  1617 => x"54738c17",
  1618 => x"23983d0d",
  1619 => x"04810b8c",
  1620 => x"17225855",
  1621 => x"fef539a8",
  1622 => x"160880c1",
  1623 => x"fc2e0981",
  1624 => x"06fee438",
  1625 => x"8c162288",
  1626 => x"80075473",
  1627 => x"8c172388",
  1628 => x"800b80cc",
  1629 => x"170cfedc",
  1630 => x"39f33d0d",
  1631 => x"7f618b11",
  1632 => x"70f8065c",
  1633 => x"55555e72",
  1634 => x"96268338",
  1635 => x"90598079",
  1636 => x"24747a26",
  1637 => x"07538054",
  1638 => x"72742e09",
  1639 => x"810680cb",
  1640 => x"387d518c",
  1641 => x"d93f7883",
  1642 => x"f72680c6",
  1643 => x"3878832a",
  1644 => x"70101010",
  1645 => x"80d4f405",
  1646 => x"8c110859",
  1647 => x"595a7678",
  1648 => x"2e83b038",
  1649 => x"841708fc",
  1650 => x"06568c17",
  1651 => x"08881808",
  1652 => x"718c120c",
  1653 => x"88120c58",
  1654 => x"75178411",
  1655 => x"08810784",
  1656 => x"120c537d",
  1657 => x"518c983f",
  1658 => x"88175473",
  1659 => x"800c8f3d",
  1660 => x"0d047889",
  1661 => x"2a79832a",
  1662 => x"5b537280",
  1663 => x"2ebf3878",
  1664 => x"862ab805",
  1665 => x"5a847327",
  1666 => x"b43880db",
  1667 => x"135a9473",
  1668 => x"27ab3878",
  1669 => x"8c2a80ee",
  1670 => x"055a80d4",
  1671 => x"73279e38",
  1672 => x"788f2a80",
  1673 => x"f7055a82",
  1674 => x"d4732791",
  1675 => x"3878922a",
  1676 => x"80fc055a",
  1677 => x"8ad47327",
  1678 => x"843880fe",
  1679 => x"5a791010",
  1680 => x"1080d4f4",
  1681 => x"058c1108",
  1682 => x"58557675",
  1683 => x"2ea33884",
  1684 => x"1708fc06",
  1685 => x"707a3155",
  1686 => x"56738f24",
  1687 => x"88d53873",
  1688 => x"8025fee6",
  1689 => x"388c1708",
  1690 => x"5776752e",
  1691 => x"098106df",
  1692 => x"38811a5a",
  1693 => x"80d58408",
  1694 => x"577680d4",
  1695 => x"fc2e82c0",
  1696 => x"38841708",
  1697 => x"fc06707a",
  1698 => x"31555673",
  1699 => x"8f2481f9",
  1700 => x"3880d4fc",
  1701 => x"0b80d588",
  1702 => x"0c80d4fc",
  1703 => x"0b80d584",
  1704 => x"0c738025",
  1705 => x"feb23883",
  1706 => x"ff762783",
  1707 => x"df387589",
  1708 => x"2a76832a",
  1709 => x"55537280",
  1710 => x"2ebf3875",
  1711 => x"862ab805",
  1712 => x"54847327",
  1713 => x"b43880db",
  1714 => x"13549473",
  1715 => x"27ab3875",
  1716 => x"8c2a80ee",
  1717 => x"055480d4",
  1718 => x"73279e38",
  1719 => x"758f2a80",
  1720 => x"f7055482",
  1721 => x"d4732791",
  1722 => x"3875922a",
  1723 => x"80fc0554",
  1724 => x"8ad47327",
  1725 => x"843880fe",
  1726 => x"54731010",
  1727 => x"1080d4f4",
  1728 => x"05881108",
  1729 => x"56587478",
  1730 => x"2e86cf38",
  1731 => x"841508fc",
  1732 => x"06537573",
  1733 => x"278d3888",
  1734 => x"15085574",
  1735 => x"782e0981",
  1736 => x"06ea388c",
  1737 => x"150880d4",
  1738 => x"f40b8405",
  1739 => x"08718c1a",
  1740 => x"0c76881a",
  1741 => x"0c788813",
  1742 => x"0c788c18",
  1743 => x"0c5d5879",
  1744 => x"53807a24",
  1745 => x"83e63872",
  1746 => x"822c8171",
  1747 => x"2b5c537a",
  1748 => x"7c268198",
  1749 => x"387b7b06",
  1750 => x"537282f1",
  1751 => x"3879fc06",
  1752 => x"84055a7a",
  1753 => x"10707d06",
  1754 => x"545b7282",
  1755 => x"e038841a",
  1756 => x"5af13988",
  1757 => x"178c1108",
  1758 => x"58587678",
  1759 => x"2e098106",
  1760 => x"fcc23882",
  1761 => x"1a5afdec",
  1762 => x"39781779",
  1763 => x"81078419",
  1764 => x"0c7080d5",
  1765 => x"880c7080",
  1766 => x"d5840c80",
  1767 => x"d4fc0b8c",
  1768 => x"120c8c11",
  1769 => x"0888120c",
  1770 => x"74810784",
  1771 => x"120c7411",
  1772 => x"75710c51",
  1773 => x"537d5188",
  1774 => x"c63f8817",
  1775 => x"54fcac39",
  1776 => x"80d4f40b",
  1777 => x"8405087a",
  1778 => x"545c7980",
  1779 => x"25fef838",
  1780 => x"82da397a",
  1781 => x"097c0670",
  1782 => x"80d4f40b",
  1783 => x"84050c5c",
  1784 => x"7a105b7a",
  1785 => x"7c268538",
  1786 => x"7a85b838",
  1787 => x"80d4f40b",
  1788 => x"88050870",
  1789 => x"841208fc",
  1790 => x"06707c31",
  1791 => x"7c72268f",
  1792 => x"72250757",
  1793 => x"575c5d55",
  1794 => x"72802e80",
  1795 => x"db38797a",
  1796 => x"1680d4ec",
  1797 => x"081b9011",
  1798 => x"5a55575b",
  1799 => x"80d4e808",
  1800 => x"ff2e8838",
  1801 => x"a08f13e0",
  1802 => x"80065776",
  1803 => x"527d5187",
  1804 => x"cf3f8008",
  1805 => x"548008ff",
  1806 => x"2e903880",
  1807 => x"08762782",
  1808 => x"99387480",
  1809 => x"d4f42e82",
  1810 => x"913880d4",
  1811 => x"f40b8805",
  1812 => x"08558415",
  1813 => x"08fc0670",
  1814 => x"7a317a72",
  1815 => x"268f7225",
  1816 => x"07525553",
  1817 => x"7283e638",
  1818 => x"74798107",
  1819 => x"84170c79",
  1820 => x"167080d4",
  1821 => x"f40b8805",
  1822 => x"0c758107",
  1823 => x"84120c54",
  1824 => x"7e525786",
  1825 => x"fa3f8817",
  1826 => x"54fae039",
  1827 => x"75832a70",
  1828 => x"54548074",
  1829 => x"24819b38",
  1830 => x"72822c81",
  1831 => x"712b80d4",
  1832 => x"f8080770",
  1833 => x"80d4f40b",
  1834 => x"84050c75",
  1835 => x"10101080",
  1836 => x"d4f40588",
  1837 => x"1108585a",
  1838 => x"5d53778c",
  1839 => x"180c7488",
  1840 => x"180c7688",
  1841 => x"190c768c",
  1842 => x"160cfcf3",
  1843 => x"39797a10",
  1844 => x"101080d4",
  1845 => x"f4057057",
  1846 => x"595d8c15",
  1847 => x"08577675",
  1848 => x"2ea33884",
  1849 => x"1708fc06",
  1850 => x"707a3155",
  1851 => x"56738f24",
  1852 => x"83ca3873",
  1853 => x"80258481",
  1854 => x"388c1708",
  1855 => x"5776752e",
  1856 => x"098106df",
  1857 => x"38881581",
  1858 => x"1b708306",
  1859 => x"555b5572",
  1860 => x"c9387c83",
  1861 => x"06537280",
  1862 => x"2efdb838",
  1863 => x"ff1df819",
  1864 => x"595d8818",
  1865 => x"08782eea",
  1866 => x"38fdb539",
  1867 => x"831a53fc",
  1868 => x"96398314",
  1869 => x"70822c81",
  1870 => x"712b80d4",
  1871 => x"f8080770",
  1872 => x"80d4f40b",
  1873 => x"84050c76",
  1874 => x"10101080",
  1875 => x"d4f40588",
  1876 => x"1108595b",
  1877 => x"5e5153fe",
  1878 => x"e13980d4",
  1879 => x"b8081758",
  1880 => x"8008762e",
  1881 => x"818d3880",
  1882 => x"d4e808ff",
  1883 => x"2e83ec38",
  1884 => x"73763118",
  1885 => x"80d4b80c",
  1886 => x"73870670",
  1887 => x"57537280",
  1888 => x"2e883888",
  1889 => x"73317015",
  1890 => x"55567614",
  1891 => x"9fff06a0",
  1892 => x"80713117",
  1893 => x"70547f53",
  1894 => x"575384e4",
  1895 => x"3f800853",
  1896 => x"8008ff2e",
  1897 => x"81a03880",
  1898 => x"d4b80816",
  1899 => x"7080d4b8",
  1900 => x"0c747580",
  1901 => x"d4f40b88",
  1902 => x"050c7476",
  1903 => x"31187081",
  1904 => x"07515556",
  1905 => x"587b80d4",
  1906 => x"f42e839c",
  1907 => x"38798f26",
  1908 => x"82cb3881",
  1909 => x"0b84150c",
  1910 => x"841508fc",
  1911 => x"06707a31",
  1912 => x"7a72268f",
  1913 => x"72250752",
  1914 => x"55537280",
  1915 => x"2efcf938",
  1916 => x"80db3980",
  1917 => x"089fff06",
  1918 => x"5372feeb",
  1919 => x"387780d4",
  1920 => x"b80c80d4",
  1921 => x"f40b8805",
  1922 => x"087b1881",
  1923 => x"0784120c",
  1924 => x"5580d4e4",
  1925 => x"08782786",
  1926 => x"387780d4",
  1927 => x"e40c80d4",
  1928 => x"e0087827",
  1929 => x"fcac3877",
  1930 => x"80d4e00c",
  1931 => x"841508fc",
  1932 => x"06707a31",
  1933 => x"7a72268f",
  1934 => x"72250752",
  1935 => x"55537280",
  1936 => x"2efca538",
  1937 => x"88398074",
  1938 => x"5456fedb",
  1939 => x"397d5183",
  1940 => x"ae3f800b",
  1941 => x"800c8f3d",
  1942 => x"0d047353",
  1943 => x"807424a9",
  1944 => x"3872822c",
  1945 => x"81712b80",
  1946 => x"d4f80807",
  1947 => x"7080d4f4",
  1948 => x"0b84050c",
  1949 => x"5d53778c",
  1950 => x"180c7488",
  1951 => x"180c7688",
  1952 => x"190c768c",
  1953 => x"160cf9b7",
  1954 => x"39831470",
  1955 => x"822c8171",
  1956 => x"2b80d4f8",
  1957 => x"08077080",
  1958 => x"d4f40b84",
  1959 => x"050c5e51",
  1960 => x"53d4397b",
  1961 => x"7b065372",
  1962 => x"fca33884",
  1963 => x"1a7b105c",
  1964 => x"5af139ff",
  1965 => x"1a811151",
  1966 => x"5af7b939",
  1967 => x"78177981",
  1968 => x"0784190c",
  1969 => x"8c180888",
  1970 => x"1908718c",
  1971 => x"120c8812",
  1972 => x"0c597080",
  1973 => x"d5880c70",
  1974 => x"80d5840c",
  1975 => x"80d4fc0b",
  1976 => x"8c120c8c",
  1977 => x"11088812",
  1978 => x"0c748107",
  1979 => x"84120c74",
  1980 => x"1175710c",
  1981 => x"5153f9bd",
  1982 => x"39751784",
  1983 => x"11088107",
  1984 => x"84120c53",
  1985 => x"8c170888",
  1986 => x"1808718c",
  1987 => x"120c8812",
  1988 => x"0c587d51",
  1989 => x"81e93f88",
  1990 => x"1754f5cf",
  1991 => x"39728415",
  1992 => x"0cf41af8",
  1993 => x"0670841e",
  1994 => x"08810607",
  1995 => x"841e0c70",
  1996 => x"1d545b85",
  1997 => x"0b84140c",
  1998 => x"850b8814",
  1999 => x"0c8f7b27",
  2000 => x"fdcf3888",
  2001 => x"1c527d51",
  2002 => x"ec9d3f80",
  2003 => x"d4f40b88",
  2004 => x"050880d4",
  2005 => x"b8085955",
  2006 => x"fdb73977",
  2007 => x"80d4b80c",
  2008 => x"7380d4e8",
  2009 => x"0cfc9139",
  2010 => x"7284150c",
  2011 => x"fda339fc",
  2012 => x"3d0d7679",
  2013 => x"71028c05",
  2014 => x"9f053357",
  2015 => x"55535583",
  2016 => x"72278a38",
  2017 => x"74830651",
  2018 => x"70802ea2",
  2019 => x"38ff1252",
  2020 => x"71ff2e93",
  2021 => x"38737370",
  2022 => x"81055534",
  2023 => x"ff125271",
  2024 => x"ff2e0981",
  2025 => x"06ef3874",
  2026 => x"800c863d",
  2027 => x"0d047474",
  2028 => x"882b7507",
  2029 => x"7071902b",
  2030 => x"07515451",
  2031 => x"8f7227a5",
  2032 => x"38727170",
  2033 => x"8405530c",
  2034 => x"72717084",
  2035 => x"05530c72",
  2036 => x"71708405",
  2037 => x"530c7271",
  2038 => x"70840553",
  2039 => x"0cf01252",
  2040 => x"718f26dd",
  2041 => x"38837227",
  2042 => x"90387271",
  2043 => x"70840553",
  2044 => x"0cfc1252",
  2045 => x"718326f2",
  2046 => x"387053ff",
  2047 => x"90390404",
  2048 => x"fd3d0d80",
  2049 => x"0b80ddb4",
  2050 => x"0c765184",
  2051 => x"ee3f8008",
  2052 => x"538008ff",
  2053 => x"2e883872",
  2054 => x"800c853d",
  2055 => x"0d0480dd",
  2056 => x"b4085473",
  2057 => x"802ef038",
  2058 => x"7574710c",
  2059 => x"5272800c",
  2060 => x"853d0d04",
  2061 => x"f93d0d79",
  2062 => x"7c557b54",
  2063 => x"8e112270",
  2064 => x"902b7090",
  2065 => x"2c555780",
  2066 => x"cdb80853",
  2067 => x"585683f3",
  2068 => x"3f800857",
  2069 => x"800b8008",
  2070 => x"24933880",
  2071 => x"d0160880",
  2072 => x"080580d0",
  2073 => x"170c7680",
  2074 => x"0c893d0d",
  2075 => x"048c1622",
  2076 => x"83dfff06",
  2077 => x"55748c17",
  2078 => x"2376800c",
  2079 => x"893d0d04",
  2080 => x"fa3d0d78",
  2081 => x"8c112270",
  2082 => x"882a7081",
  2083 => x"06515758",
  2084 => x"5674a938",
  2085 => x"8c162283",
  2086 => x"dfff0655",
  2087 => x"748c1723",
  2088 => x"7a547953",
  2089 => x"8e162270",
  2090 => x"902b7090",
  2091 => x"2c545680",
  2092 => x"cdb80852",
  2093 => x"5681b23f",
  2094 => x"883d0d04",
  2095 => x"82548053",
  2096 => x"8e162270",
  2097 => x"902b7090",
  2098 => x"2c545680",
  2099 => x"cdb80852",
  2100 => x"5782b83f",
  2101 => x"8c162283",
  2102 => x"dfff0655",
  2103 => x"748c1723",
  2104 => x"7a547953",
  2105 => x"8e162270",
  2106 => x"902b7090",
  2107 => x"2c545680",
  2108 => x"cdb80852",
  2109 => x"5680f23f",
  2110 => x"883d0d04",
  2111 => x"f93d0d79",
  2112 => x"7c557b54",
  2113 => x"8e112270",
  2114 => x"902b7090",
  2115 => x"2c555780",
  2116 => x"cdb80853",
  2117 => x"585681f3",
  2118 => x"3f800857",
  2119 => x"8008ff2e",
  2120 => x"99388c16",
  2121 => x"22a08007",
  2122 => x"55748c17",
  2123 => x"23800880",
  2124 => x"d0170c76",
  2125 => x"800c893d",
  2126 => x"0d048c16",
  2127 => x"2283dfff",
  2128 => x"0655748c",
  2129 => x"17237680",
  2130 => x"0c893d0d",
  2131 => x"04fe3d0d",
  2132 => x"748e1122",
  2133 => x"70902b70",
  2134 => x"902c5551",
  2135 => x"515380cd",
  2136 => x"b80851bd",
  2137 => x"3f843d0d",
  2138 => x"04fb3d0d",
  2139 => x"800b80dd",
  2140 => x"b40c7a53",
  2141 => x"79527851",
  2142 => x"82fc3f80",
  2143 => x"08558008",
  2144 => x"ff2e8838",
  2145 => x"74800c87",
  2146 => x"3d0d0480",
  2147 => x"ddb40856",
  2148 => x"75802ef0",
  2149 => x"38777671",
  2150 => x"0c547480",
  2151 => x"0c873d0d",
  2152 => x"04fd3d0d",
  2153 => x"800b80dd",
  2154 => x"b40c7651",
  2155 => x"84c63f80",
  2156 => x"08538008",
  2157 => x"ff2e8838",
  2158 => x"72800c85",
  2159 => x"3d0d0480",
  2160 => x"ddb40854",
  2161 => x"73802ef0",
  2162 => x"38757471",
  2163 => x"0c527280",
  2164 => x"0c853d0d",
  2165 => x"04fc3d0d",
  2166 => x"800b80dd",
  2167 => x"b40c7852",
  2168 => x"775186ac",
  2169 => x"3f800854",
  2170 => x"8008ff2e",
  2171 => x"88387380",
  2172 => x"0c863d0d",
  2173 => x"0480ddb4",
  2174 => x"08557480",
  2175 => x"2ef03876",
  2176 => x"75710c53",
  2177 => x"73800c86",
  2178 => x"3d0d04fb",
  2179 => x"3d0d800b",
  2180 => x"80ddb40c",
  2181 => x"7a537952",
  2182 => x"78518489",
  2183 => x"3f800855",
  2184 => x"8008ff2e",
  2185 => x"88387480",
  2186 => x"0c873d0d",
  2187 => x"0480ddb4",
  2188 => x"08567580",
  2189 => x"2ef03877",
  2190 => x"76710c54",
  2191 => x"74800c87",
  2192 => x"3d0d04fb",
  2193 => x"3d0d800b",
  2194 => x"80ddb40c",
  2195 => x"7a537952",
  2196 => x"78518296",
  2197 => x"3f800855",
  2198 => x"8008ff2e",
  2199 => x"88387480",
  2200 => x"0c873d0d",
  2201 => x"0480ddb4",
  2202 => x"08567580",
  2203 => x"2ef03877",
  2204 => x"76710c54",
  2205 => x"74800c87",
  2206 => x"3d0d04fe",
  2207 => x"3d0d80dd",
  2208 => x"a4085170",
  2209 => x"8a3880dd",
  2210 => x"b87080dd",
  2211 => x"a40c5170",
  2212 => x"75125252",
  2213 => x"ff537087",
  2214 => x"fb808026",
  2215 => x"88387080",
  2216 => x"dda40c71",
  2217 => x"5372800c",
  2218 => x"843d0d04",
  2219 => x"fd3d0d80",
  2220 => x"0b80cdac",
  2221 => x"08545472",
  2222 => x"812e9b38",
  2223 => x"7380dda8",
  2224 => x"0cc3e33f",
  2225 => x"c2ba3f80",
  2226 => x"dcfc5281",
  2227 => x"51c5a93f",
  2228 => x"80085185",
  2229 => x"bb3f7280",
  2230 => x"dda80cc3",
  2231 => x"c93fc2a0",
  2232 => x"3f80dcfc",
  2233 => x"528151c5",
  2234 => x"8f3f8008",
  2235 => x"5185a13f",
  2236 => x"00ff3900",
  2237 => x"ff39f53d",
  2238 => x"0d7e6080",
  2239 => x"dda80870",
  2240 => x"5b585b5b",
  2241 => x"7580c238",
  2242 => x"777a25a1",
  2243 => x"38771b70",
  2244 => x"337081ff",
  2245 => x"06585859",
  2246 => x"758a2e98",
  2247 => x"387681ff",
  2248 => x"0651c2e1",
  2249 => x"3f811858",
  2250 => x"797824e1",
  2251 => x"3879800c",
  2252 => x"8d3d0d04",
  2253 => x"8d51c2cd",
  2254 => x"3f783370",
  2255 => x"81ff0652",
  2256 => x"57c2c23f",
  2257 => x"811858e0",
  2258 => x"3979557a",
  2259 => x"547d5385",
  2260 => x"528d3dfc",
  2261 => x"0551c1ea",
  2262 => x"3f800856",
  2263 => x"84ab3f7b",
  2264 => x"80080c75",
  2265 => x"800c8d3d",
  2266 => x"0d04f63d",
  2267 => x"0d7d7f80",
  2268 => x"dda80870",
  2269 => x"5b585a5a",
  2270 => x"7580c138",
  2271 => x"777925b3",
  2272 => x"38c1dd3f",
  2273 => x"800881ff",
  2274 => x"06708d32",
  2275 => x"7030709f",
  2276 => x"2a515157",
  2277 => x"57768a2e",
  2278 => x"80c33875",
  2279 => x"802ebe38",
  2280 => x"771a5676",
  2281 => x"76347651",
  2282 => x"c1db3f81",
  2283 => x"18587878",
  2284 => x"24cf3877",
  2285 => x"5675800c",
  2286 => x"8c3d0d04",
  2287 => x"78557954",
  2288 => x"7c538452",
  2289 => x"8c3dfc05",
  2290 => x"51c0f73f",
  2291 => x"80085683",
  2292 => x"b83f7a80",
  2293 => x"080c7580",
  2294 => x"0c8c3d0d",
  2295 => x"04771a56",
  2296 => x"8a763481",
  2297 => x"18588d51",
  2298 => x"c19b3f8a",
  2299 => x"51c1963f",
  2300 => x"7756c239",
  2301 => x"fb3d0d80",
  2302 => x"dda80870",
  2303 => x"56547388",
  2304 => x"3874800c",
  2305 => x"873d0d04",
  2306 => x"77538352",
  2307 => x"873dfc05",
  2308 => x"51c0af3f",
  2309 => x"80085482",
  2310 => x"f03f7580",
  2311 => x"080c7380",
  2312 => x"0c873d0d",
  2313 => x"04fa3d0d",
  2314 => x"80dda808",
  2315 => x"802ea238",
  2316 => x"7a557954",
  2317 => x"78538652",
  2318 => x"883dfc05",
  2319 => x"51c0833f",
  2320 => x"80085682",
  2321 => x"c43f7680",
  2322 => x"080c7580",
  2323 => x"0c883d0d",
  2324 => x"0482b63f",
  2325 => x"9d0b8008",
  2326 => x"0cff0b80",
  2327 => x"0c883d0d",
  2328 => x"04fb3d0d",
  2329 => x"77795656",
  2330 => x"80705454",
  2331 => x"7375259f",
  2332 => x"38741010",
  2333 => x"10f80552",
  2334 => x"72167033",
  2335 => x"70742b76",
  2336 => x"078116f8",
  2337 => x"16565656",
  2338 => x"51517473",
  2339 => x"24ea3873",
  2340 => x"800c873d",
  2341 => x"0d04fc3d",
  2342 => x"0d767855",
  2343 => x"55bc5380",
  2344 => x"527351f5",
  2345 => x"ca3f8452",
  2346 => x"7451ffb5",
  2347 => x"3f800874",
  2348 => x"23845284",
  2349 => x"1551ffa9",
  2350 => x"3f800882",
  2351 => x"15238452",
  2352 => x"881551ff",
  2353 => x"9c3f8008",
  2354 => x"84150c84",
  2355 => x"528c1551",
  2356 => x"ff8f3f80",
  2357 => x"08881523",
  2358 => x"84529015",
  2359 => x"51ff823f",
  2360 => x"80088a15",
  2361 => x"23845294",
  2362 => x"1551fef5",
  2363 => x"3f80088c",
  2364 => x"15238452",
  2365 => x"981551fe",
  2366 => x"e83f8008",
  2367 => x"8e152388",
  2368 => x"529c1551",
  2369 => x"fedb3f80",
  2370 => x"0890150c",
  2371 => x"863d0d04",
  2372 => x"e93d0d6a",
  2373 => x"80dda808",
  2374 => x"57577593",
  2375 => x"3880c080",
  2376 => x"0b84180c",
  2377 => x"75ac180c",
  2378 => x"75800c99",
  2379 => x"3d0d0489",
  2380 => x"3d70556a",
  2381 => x"54558a52",
  2382 => x"993dffbc",
  2383 => x"0551ffbe",
  2384 => x"813f8008",
  2385 => x"77537552",
  2386 => x"56fecb3f",
  2387 => x"bc3f7780",
  2388 => x"080c7580",
  2389 => x"0c993d0d",
  2390 => x"04fc3d0d",
  2391 => x"815480dd",
  2392 => x"a8088838",
  2393 => x"73800c86",
  2394 => x"3d0d0476",
  2395 => x"5397b952",
  2396 => x"863dfc05",
  2397 => x"51ffbdca",
  2398 => x"3f800854",
  2399 => x"8c3f7480",
  2400 => x"080c7380",
  2401 => x"0c863d0d",
  2402 => x"0480cdb8",
  2403 => x"08800c04",
  2404 => x"f73d0d7b",
  2405 => x"80cdb808",
  2406 => x"82c81108",
  2407 => x"5a545a77",
  2408 => x"802e80da",
  2409 => x"38818818",
  2410 => x"841908ff",
  2411 => x"0581712b",
  2412 => x"59555980",
  2413 => x"742480ea",
  2414 => x"38807424",
  2415 => x"b5387382",
  2416 => x"2b781188",
  2417 => x"05565681",
  2418 => x"80190877",
  2419 => x"06537280",
  2420 => x"2eb63878",
  2421 => x"16700853",
  2422 => x"53795174",
  2423 => x"0853722d",
  2424 => x"ff14fc17",
  2425 => x"fc177981",
  2426 => x"2c5a5757",
  2427 => x"54738025",
  2428 => x"d6387708",
  2429 => x"5877ffad",
  2430 => x"3880cdb8",
  2431 => x"0853bc13",
  2432 => x"08a53879",
  2433 => x"51f9e93f",
  2434 => x"74085372",
  2435 => x"2dff14fc",
  2436 => x"17fc1779",
  2437 => x"812c5a57",
  2438 => x"57547380",
  2439 => x"25ffa838",
  2440 => x"d1398057",
  2441 => x"ff933972",
  2442 => x"51bc1308",
  2443 => x"53722d79",
  2444 => x"51f9bd3f",
  2445 => x"ff3d0d80",
  2446 => x"dd840bfc",
  2447 => x"05700852",
  2448 => x"5270ff2e",
  2449 => x"9138702d",
  2450 => x"fc127008",
  2451 => x"525270ff",
  2452 => x"2e098106",
  2453 => x"f138833d",
  2454 => x"0d0404ff",
  2455 => x"bdb53f04",
  2456 => x"00000040",
  2457 => x"48656c6c",
  2458 => x"6f20776f",
  2459 => x"726c6420",
  2460 => x"310a0000",
  2461 => x"48656c6c",
  2462 => x"6f20776f",
  2463 => x"726c6420",
  2464 => x"320a0000",
  2465 => x"0a000000",
  2466 => x"43000000",
  2467 => x"64756d6d",
  2468 => x"792e6578",
  2469 => x"65000000",
  2470 => x"00ffffff",
  2471 => x"ff00ffff",
  2472 => x"ffff00ff",
  2473 => x"ffffff00",
  2474 => x"00000000",
  2475 => x"00000000",
  2476 => x"00000000",
  2477 => x"00002e8c",
  2478 => x"000026bc",
  2479 => x"00000000",
  2480 => x"00002924",
  2481 => x"00002980",
  2482 => x"000029dc",
  2483 => x"00000000",
  2484 => x"00000000",
  2485 => x"00000000",
  2486 => x"00000000",
  2487 => x"00000000",
  2488 => x"00000000",
  2489 => x"00000000",
  2490 => x"00000000",
  2491 => x"00000000",
  2492 => x"00002688",
  2493 => x"00000000",
  2494 => x"00000000",
  2495 => x"00000000",
  2496 => x"00000000",
  2497 => x"00000000",
  2498 => x"00000000",
  2499 => x"00000000",
  2500 => x"00000000",
  2501 => x"00000000",
  2502 => x"00000000",
  2503 => x"00000000",
  2504 => x"00000000",
  2505 => x"00000000",
  2506 => x"00000000",
  2507 => x"00000000",
  2508 => x"00000000",
  2509 => x"00000000",
  2510 => x"00000000",
  2511 => x"00000000",
  2512 => x"00000000",
  2513 => x"00000000",
  2514 => x"00000000",
  2515 => x"00000000",
  2516 => x"00000000",
  2517 => x"00000000",
  2518 => x"00000000",
  2519 => x"00000000",
  2520 => x"00000000",
  2521 => x"00000001",
  2522 => x"330eabcd",
  2523 => x"1234e66d",
  2524 => x"deec0005",
  2525 => x"000b0000",
  2526 => x"00000000",
  2527 => x"00000000",
  2528 => x"00000000",
  2529 => x"00000000",
  2530 => x"00000000",
  2531 => x"00000000",
  2532 => x"00000000",
  2533 => x"00000000",
  2534 => x"00000000",
  2535 => x"00000000",
  2536 => x"00000000",
  2537 => x"00000000",
  2538 => x"00000000",
  2539 => x"00000000",
  2540 => x"00000000",
  2541 => x"00000000",
  2542 => x"00000000",
  2543 => x"00000000",
  2544 => x"00000000",
  2545 => x"00000000",
  2546 => x"00000000",
  2547 => x"00000000",
  2548 => x"00000000",
  2549 => x"00000000",
  2550 => x"00000000",
  2551 => x"00000000",
  2552 => x"00000000",
  2553 => x"00000000",
  2554 => x"00000000",
  2555 => x"00000000",
  2556 => x"00000000",
  2557 => x"00000000",
  2558 => x"00000000",
  2559 => x"00000000",
  2560 => x"00000000",
  2561 => x"00000000",
  2562 => x"00000000",
  2563 => x"00000000",
  2564 => x"00000000",
  2565 => x"00000000",
  2566 => x"00000000",
  2567 => x"00000000",
  2568 => x"00000000",
  2569 => x"00000000",
  2570 => x"00000000",
  2571 => x"00000000",
  2572 => x"00000000",
  2573 => x"00000000",
  2574 => x"00000000",
  2575 => x"00000000",
  2576 => x"00000000",
  2577 => x"00000000",
  2578 => x"00000000",
  2579 => x"00000000",
  2580 => x"00000000",
  2581 => x"00000000",
  2582 => x"00000000",
  2583 => x"00000000",
  2584 => x"00000000",
  2585 => x"00000000",
  2586 => x"00000000",
  2587 => x"00000000",
  2588 => x"00000000",
  2589 => x"00000000",
  2590 => x"00000000",
  2591 => x"00000000",
  2592 => x"00000000",
  2593 => x"00000000",
  2594 => x"00000000",
  2595 => x"00000000",
  2596 => x"00000000",
  2597 => x"00000000",
  2598 => x"00000000",
  2599 => x"00000000",
  2600 => x"00000000",
  2601 => x"00000000",
  2602 => x"00000000",
  2603 => x"00000000",
  2604 => x"00000000",
  2605 => x"00000000",
  2606 => x"00000000",
  2607 => x"00000000",
  2608 => x"00000000",
  2609 => x"00000000",
  2610 => x"00000000",
  2611 => x"00000000",
  2612 => x"00000000",
  2613 => x"00000000",
  2614 => x"00000000",
  2615 => x"00000000",
  2616 => x"00000000",
  2617 => x"00000000",
  2618 => x"00000000",
  2619 => x"00000000",
  2620 => x"00000000",
  2621 => x"00000000",
  2622 => x"00000000",
  2623 => x"00000000",
  2624 => x"00000000",
  2625 => x"00000000",
  2626 => x"00000000",
  2627 => x"00000000",
  2628 => x"00000000",
  2629 => x"00000000",
  2630 => x"00000000",
  2631 => x"00000000",
  2632 => x"00000000",
  2633 => x"00000000",
  2634 => x"00000000",
  2635 => x"00000000",
  2636 => x"00000000",
  2637 => x"00000000",
  2638 => x"00000000",
  2639 => x"00000000",
  2640 => x"00000000",
  2641 => x"00000000",
  2642 => x"00000000",
  2643 => x"00000000",
  2644 => x"00000000",
  2645 => x"00000000",
  2646 => x"00000000",
  2647 => x"00000000",
  2648 => x"00000000",
  2649 => x"00000000",
  2650 => x"00000000",
  2651 => x"00000000",
  2652 => x"00000000",
  2653 => x"00000000",
  2654 => x"00000000",
  2655 => x"00000000",
  2656 => x"00000000",
  2657 => x"00000000",
  2658 => x"00000000",
  2659 => x"00000000",
  2660 => x"00000000",
  2661 => x"00000000",
  2662 => x"00000000",
  2663 => x"00000000",
  2664 => x"00000000",
  2665 => x"00000000",
  2666 => x"00000000",
  2667 => x"00000000",
  2668 => x"00000000",
  2669 => x"00000000",
  2670 => x"00000000",
  2671 => x"00000000",
  2672 => x"00000000",
  2673 => x"00000000",
  2674 => x"00000000",
  2675 => x"00000000",
  2676 => x"00000000",
  2677 => x"00000000",
  2678 => x"00000000",
  2679 => x"00000000",
  2680 => x"00000000",
  2681 => x"00000000",
  2682 => x"00000000",
  2683 => x"00000000",
  2684 => x"00000000",
  2685 => x"00000000",
  2686 => x"00000000",
  2687 => x"00000000",
  2688 => x"00000000",
  2689 => x"00000000",
  2690 => x"00000000",
  2691 => x"00000000",
  2692 => x"00000000",
  2693 => x"00000000",
  2694 => x"00000000",
  2695 => x"00000000",
  2696 => x"00000000",
  2697 => x"00000000",
  2698 => x"00000000",
  2699 => x"00000000",
  2700 => x"00000000",
  2701 => x"00000000",
  2702 => x"00000000",
  2703 => x"00000000",
  2704 => x"00000000",
  2705 => x"00000000",
  2706 => x"00000000",
  2707 => x"00000000",
  2708 => x"00000000",
  2709 => x"00000000",
  2710 => x"00000000",
  2711 => x"00000000",
  2712 => x"00000000",
  2713 => x"00000000",
  2714 => x"ffffffff",
  2715 => x"00000000",
  2716 => x"00020000",
  2717 => x"00000000",
  2718 => x"00000000",
  2719 => x"00002a74",
  2720 => x"00002a74",
  2721 => x"00002a7c",
  2722 => x"00002a7c",
  2723 => x"00002a84",
  2724 => x"00002a84",
  2725 => x"00002a8c",
  2726 => x"00002a8c",
  2727 => x"00002a94",
  2728 => x"00002a94",
  2729 => x"00002a9c",
  2730 => x"00002a9c",
  2731 => x"00002aa4",
  2732 => x"00002aa4",
  2733 => x"00002aac",
  2734 => x"00002aac",
  2735 => x"00002ab4",
  2736 => x"00002ab4",
  2737 => x"00002abc",
  2738 => x"00002abc",
  2739 => x"00002ac4",
  2740 => x"00002ac4",
  2741 => x"00002acc",
  2742 => x"00002acc",
  2743 => x"00002ad4",
  2744 => x"00002ad4",
  2745 => x"00002adc",
  2746 => x"00002adc",
  2747 => x"00002ae4",
  2748 => x"00002ae4",
  2749 => x"00002aec",
  2750 => x"00002aec",
  2751 => x"00002af4",
  2752 => x"00002af4",
  2753 => x"00002afc",
  2754 => x"00002afc",
  2755 => x"00002b04",
  2756 => x"00002b04",
  2757 => x"00002b0c",
  2758 => x"00002b0c",
  2759 => x"00002b14",
  2760 => x"00002b14",
  2761 => x"00002b1c",
  2762 => x"00002b1c",
  2763 => x"00002b24",
  2764 => x"00002b24",
  2765 => x"00002b2c",
  2766 => x"00002b2c",
  2767 => x"00002b34",
  2768 => x"00002b34",
  2769 => x"00002b3c",
  2770 => x"00002b3c",
  2771 => x"00002b44",
  2772 => x"00002b44",
  2773 => x"00002b4c",
  2774 => x"00002b4c",
  2775 => x"00002b54",
  2776 => x"00002b54",
  2777 => x"00002b5c",
  2778 => x"00002b5c",
  2779 => x"00002b64",
  2780 => x"00002b64",
  2781 => x"00002b6c",
  2782 => x"00002b6c",
  2783 => x"00002b74",
  2784 => x"00002b74",
  2785 => x"00002b7c",
  2786 => x"00002b7c",
  2787 => x"00002b84",
  2788 => x"00002b84",
  2789 => x"00002b8c",
  2790 => x"00002b8c",
  2791 => x"00002b94",
  2792 => x"00002b94",
  2793 => x"00002b9c",
  2794 => x"00002b9c",
  2795 => x"00002ba4",
  2796 => x"00002ba4",
  2797 => x"00002bac",
  2798 => x"00002bac",
  2799 => x"00002bb4",
  2800 => x"00002bb4",
  2801 => x"00002bbc",
  2802 => x"00002bbc",
  2803 => x"00002bc4",
  2804 => x"00002bc4",
  2805 => x"00002bcc",
  2806 => x"00002bcc",
  2807 => x"00002bd4",
  2808 => x"00002bd4",
  2809 => x"00002bdc",
  2810 => x"00002bdc",
  2811 => x"00002be4",
  2812 => x"00002be4",
  2813 => x"00002bec",
  2814 => x"00002bec",
  2815 => x"00002bf4",
  2816 => x"00002bf4",
  2817 => x"00002bfc",
  2818 => x"00002bfc",
  2819 => x"00002c04",
  2820 => x"00002c04",
  2821 => x"00002c0c",
  2822 => x"00002c0c",
  2823 => x"00002c14",
  2824 => x"00002c14",
  2825 => x"00002c1c",
  2826 => x"00002c1c",
  2827 => x"00002c24",
  2828 => x"00002c24",
  2829 => x"00002c2c",
  2830 => x"00002c2c",
  2831 => x"00002c34",
  2832 => x"00002c34",
  2833 => x"00002c3c",
  2834 => x"00002c3c",
  2835 => x"00002c44",
  2836 => x"00002c44",
  2837 => x"00002c4c",
  2838 => x"00002c4c",
  2839 => x"00002c54",
  2840 => x"00002c54",
  2841 => x"00002c5c",
  2842 => x"00002c5c",
  2843 => x"00002c64",
  2844 => x"00002c64",
  2845 => x"00002c6c",
  2846 => x"00002c6c",
  2847 => x"00002c74",
  2848 => x"00002c74",
  2849 => x"00002c7c",
  2850 => x"00002c7c",
  2851 => x"00002c84",
  2852 => x"00002c84",
  2853 => x"00002c8c",
  2854 => x"00002c8c",
  2855 => x"00002c94",
  2856 => x"00002c94",
  2857 => x"00002c9c",
  2858 => x"00002c9c",
  2859 => x"00002ca4",
  2860 => x"00002ca4",
  2861 => x"00002cac",
  2862 => x"00002cac",
  2863 => x"00002cb4",
  2864 => x"00002cb4",
  2865 => x"00002cbc",
  2866 => x"00002cbc",
  2867 => x"00002cc4",
  2868 => x"00002cc4",
  2869 => x"00002ccc",
  2870 => x"00002ccc",
  2871 => x"00002cd4",
  2872 => x"00002cd4",
  2873 => x"00002cdc",
  2874 => x"00002cdc",
  2875 => x"00002ce4",
  2876 => x"00002ce4",
  2877 => x"00002cec",
  2878 => x"00002cec",
  2879 => x"00002cf4",
  2880 => x"00002cf4",
  2881 => x"00002cfc",
  2882 => x"00002cfc",
  2883 => x"00002d04",
  2884 => x"00002d04",
  2885 => x"00002d0c",
  2886 => x"00002d0c",
  2887 => x"00002d14",
  2888 => x"00002d14",
  2889 => x"00002d1c",
  2890 => x"00002d1c",
  2891 => x"00002d24",
  2892 => x"00002d24",
  2893 => x"00002d2c",
  2894 => x"00002d2c",
  2895 => x"00002d34",
  2896 => x"00002d34",
  2897 => x"00002d3c",
  2898 => x"00002d3c",
  2899 => x"00002d44",
  2900 => x"00002d44",
  2901 => x"00002d4c",
  2902 => x"00002d4c",
  2903 => x"00002d54",
  2904 => x"00002d54",
  2905 => x"00002d5c",
  2906 => x"00002d5c",
  2907 => x"00002d64",
  2908 => x"00002d64",
  2909 => x"00002d6c",
  2910 => x"00002d6c",
  2911 => x"00002d74",
  2912 => x"00002d74",
  2913 => x"00002d7c",
  2914 => x"00002d7c",
  2915 => x"00002d84",
  2916 => x"00002d84",
  2917 => x"00002d8c",
  2918 => x"00002d8c",
  2919 => x"00002d94",
  2920 => x"00002d94",
  2921 => x"00002d9c",
  2922 => x"00002d9c",
  2923 => x"00002da4",
  2924 => x"00002da4",
  2925 => x"00002dac",
  2926 => x"00002dac",
  2927 => x"00002db4",
  2928 => x"00002db4",
  2929 => x"00002dbc",
  2930 => x"00002dbc",
  2931 => x"00002dc4",
  2932 => x"00002dc4",
  2933 => x"00002dcc",
  2934 => x"00002dcc",
  2935 => x"00002dd4",
  2936 => x"00002dd4",
  2937 => x"00002ddc",
  2938 => x"00002ddc",
  2939 => x"00002de4",
  2940 => x"00002de4",
  2941 => x"00002dec",
  2942 => x"00002dec",
  2943 => x"00002df4",
  2944 => x"00002df4",
  2945 => x"00002dfc",
  2946 => x"00002dfc",
  2947 => x"00002e04",
  2948 => x"00002e04",
  2949 => x"00002e0c",
  2950 => x"00002e0c",
  2951 => x"00002e14",
  2952 => x"00002e14",
  2953 => x"00002e1c",
  2954 => x"00002e1c",
  2955 => x"00002e24",
  2956 => x"00002e24",
  2957 => x"00002e2c",
  2958 => x"00002e2c",
  2959 => x"00002e34",
  2960 => x"00002e34",
  2961 => x"00002e3c",
  2962 => x"00002e3c",
  2963 => x"00002e44",
  2964 => x"00002e44",
  2965 => x"00002e4c",
  2966 => x"00002e4c",
  2967 => x"00002e54",
  2968 => x"00002e54",
  2969 => x"00002e5c",
  2970 => x"00002e5c",
  2971 => x"00002e64",
  2972 => x"00002e64",
  2973 => x"00002e6c",
  2974 => x"00002e6c",
  2975 => x"0000268c",
  2976 => x"ffffffff",
  2977 => x"00000000",
  2978 => x"ffffffff",
  2979 => x"00000000",
  2980 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
