-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"0b91a00c",
     3 => x"3a0b0b0b",
     4 => x"8ee80400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"0b8fa82d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0b91",
   162 => x"8c738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0b8a",
   171 => x"ec2d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0b8c",
   179 => x"9e2d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"0b919c0c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"81f33f88",
   257 => x"c83f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"53510491",
   280 => x"9c08802e",
   281 => x"a13891a0",
   282 => x"08822eb9",
   283 => x"38838080",
   284 => x"0b0b0b0b",
   285 => x"98cc0c82",
   286 => x"a0800b98",
   287 => x"d00c8290",
   288 => x"800b98d4",
   289 => x"0c04f880",
   290 => x"8080a40b",
   291 => x"0b0b0b98",
   292 => x"cc0cf880",
   293 => x"8082800b",
   294 => x"98d00cf8",
   295 => x"80808480",
   296 => x"0b98d40c",
   297 => x"0480c0a8",
   298 => x"808c0b0b",
   299 => x"0b0b98cc",
   300 => x"0c80c0a8",
   301 => x"80940b98",
   302 => x"d00c0b0b",
   303 => x"0b90f80b",
   304 => x"98d40c04",
   305 => x"ff3d0d98",
   306 => x"d8335170",
   307 => x"a33891a8",
   308 => x"08700852",
   309 => x"5270802e",
   310 => x"92388412",
   311 => x"91a80c70",
   312 => x"2d91a808",
   313 => x"70085252",
   314 => x"70f03881",
   315 => x"0b98d834",
   316 => x"833d0d04",
   317 => x"04803d0d",
   318 => x"0b0b0b98",
   319 => x"c808802e",
   320 => x"8e380b0b",
   321 => x"0b0b800b",
   322 => x"802e0981",
   323 => x"06853882",
   324 => x"3d0d040b",
   325 => x"0b0b98c8",
   326 => x"510b0b0b",
   327 => x"f5e23f82",
   328 => x"3d0d0404",
   329 => x"fe3d0d80",
   330 => x"0b91ac08",
   331 => x"71710c52",
   332 => x"91b00852",
   333 => x"5381710c",
   334 => x"81732b81",
   335 => x"1491b008",
   336 => x"5354710c",
   337 => x"72883270",
   338 => x"30707207",
   339 => x"9f2c7506",
   340 => x"55525280",
   341 => x"528386cf",
   342 => x"51ce1151",
   343 => x"708025f9",
   344 => x"38811252",
   345 => x"81c77227",
   346 => x"ec38cd39",
   347 => x"8c08028c",
   348 => x"0cf93d0d",
   349 => x"800b8c08",
   350 => x"fc050c8c",
   351 => x"08880508",
   352 => x"8025ab38",
   353 => x"8c088805",
   354 => x"08308c08",
   355 => x"88050c80",
   356 => x"0b8c08f4",
   357 => x"050c8c08",
   358 => x"fc050888",
   359 => x"38810b8c",
   360 => x"08f4050c",
   361 => x"8c08f405",
   362 => x"088c08fc",
   363 => x"050c8c08",
   364 => x"8c050880",
   365 => x"25ab388c",
   366 => x"088c0508",
   367 => x"308c088c",
   368 => x"050c800b",
   369 => x"8c08f005",
   370 => x"0c8c08fc",
   371 => x"05088838",
   372 => x"810b8c08",
   373 => x"f0050c8c",
   374 => x"08f00508",
   375 => x"8c08fc05",
   376 => x"0c80538c",
   377 => x"088c0508",
   378 => x"528c0888",
   379 => x"05085181",
   380 => x"a73f8008",
   381 => x"708c08f8",
   382 => x"050c548c",
   383 => x"08fc0508",
   384 => x"802e8c38",
   385 => x"8c08f805",
   386 => x"08308c08",
   387 => x"f8050c8c",
   388 => x"08f80508",
   389 => x"70800c54",
   390 => x"893d0d8c",
   391 => x"0c048c08",
   392 => x"028c0cfb",
   393 => x"3d0d800b",
   394 => x"8c08fc05",
   395 => x"0c8c0888",
   396 => x"05088025",
   397 => x"93388c08",
   398 => x"88050830",
   399 => x"8c088805",
   400 => x"0c810b8c",
   401 => x"08fc050c",
   402 => x"8c088c05",
   403 => x"0880258c",
   404 => x"388c088c",
   405 => x"0508308c",
   406 => x"088c050c",
   407 => x"81538c08",
   408 => x"8c050852",
   409 => x"8c088805",
   410 => x"0851ad3f",
   411 => x"8008708c",
   412 => x"08f8050c",
   413 => x"548c08fc",
   414 => x"0508802e",
   415 => x"8c388c08",
   416 => x"f8050830",
   417 => x"8c08f805",
   418 => x"0c8c08f8",
   419 => x"05087080",
   420 => x"0c54873d",
   421 => x"0d8c0c04",
   422 => x"8c08028c",
   423 => x"0cfd3d0d",
   424 => x"810b8c08",
   425 => x"fc050c80",
   426 => x"0b8c08f8",
   427 => x"050c8c08",
   428 => x"8c05088c",
   429 => x"08880508",
   430 => x"27ac388c",
   431 => x"08fc0508",
   432 => x"802ea338",
   433 => x"800b8c08",
   434 => x"8c050824",
   435 => x"99388c08",
   436 => x"8c050810",
   437 => x"8c088c05",
   438 => x"0c8c08fc",
   439 => x"0508108c",
   440 => x"08fc050c",
   441 => x"c9398c08",
   442 => x"fc050880",
   443 => x"2e80c938",
   444 => x"8c088c05",
   445 => x"088c0888",
   446 => x"050826a1",
   447 => x"388c0888",
   448 => x"05088c08",
   449 => x"8c050831",
   450 => x"8c088805",
   451 => x"0c8c08f8",
   452 => x"05088c08",
   453 => x"fc050807",
   454 => x"8c08f805",
   455 => x"0c8c08fc",
   456 => x"0508812a",
   457 => x"8c08fc05",
   458 => x"0c8c088c",
   459 => x"0508812a",
   460 => x"8c088c05",
   461 => x"0cffaf39",
   462 => x"8c089005",
   463 => x"08802e8f",
   464 => x"388c0888",
   465 => x"0508708c",
   466 => x"08f4050c",
   467 => x"518d398c",
   468 => x"08f80508",
   469 => x"708c08f4",
   470 => x"050c518c",
   471 => x"08f40508",
   472 => x"800c853d",
   473 => x"0d8c0c04",
   474 => x"fd3d0d80",
   475 => x"0b91a008",
   476 => x"54547281",
   477 => x"2e983873",
   478 => x"98dc0cf9",
   479 => x"e23ff980",
   480 => x"3f91b452",
   481 => x"8151fb9c",
   482 => x"3f800851",
   483 => x"9e3f7298",
   484 => x"dc0cf9cb",
   485 => x"3ff8e93f",
   486 => x"91b45281",
   487 => x"51fb853f",
   488 => x"80085187",
   489 => x"3f00ff39",
   490 => x"00ff39f7",
   491 => x"3d0d7b91",
   492 => x"b80882c8",
   493 => x"11085a54",
   494 => x"5a77802e",
   495 => x"80d93881",
   496 => x"88188419",
   497 => x"08ff0581",
   498 => x"712b5955",
   499 => x"59807424",
   500 => x"80e93880",
   501 => x"7424b538",
   502 => x"73822b78",
   503 => x"11880556",
   504 => x"56818019",
   505 => x"08770653",
   506 => x"72802eb5",
   507 => x"38781670",
   508 => x"08535379",
   509 => x"51740853",
   510 => x"722dff14",
   511 => x"fc17fc17",
   512 => x"79812c5a",
   513 => x"57575473",
   514 => x"8025d638",
   515 => x"77085877",
   516 => x"ffad3891",
   517 => x"b80853bc",
   518 => x"1308a538",
   519 => x"7951ff85",
   520 => x"3f740853",
   521 => x"722dff14",
   522 => x"fc17fc17",
   523 => x"79812c5a",
   524 => x"57575473",
   525 => x"8025ffa9",
   526 => x"38d23980",
   527 => x"57ff9439",
   528 => x"7251bc13",
   529 => x"0853722d",
   530 => x"7951fed9",
   531 => x"3fff3d0d",
   532 => x"98bc0bfc",
   533 => x"05700852",
   534 => x"5270ff2e",
   535 => x"9138702d",
   536 => x"fc127008",
   537 => x"525270ff",
   538 => x"2e098106",
   539 => x"f138833d",
   540 => x"0d0404f8",
   541 => x"cf3f0400",
   542 => x"00000040",
   543 => x"64756d6d",
   544 => x"792e6578",
   545 => x"65000000",
   546 => x"43000000",
   547 => x"00ffffff",
   548 => x"ff00ffff",
   549 => x"ffff00ff",
   550 => x"ffffff00",
   551 => x"00000000",
   552 => x"00000000",
   553 => x"00000000",
   554 => x"00000c44",
   555 => x"0c000004",
   556 => x"0c000000",
   557 => x"0000087c",
   558 => x"000008bc",
   559 => x"00000000",
   560 => x"00000b24",
   561 => x"00000b80",
   562 => x"00000bdc",
   563 => x"00000000",
   564 => x"00000000",
   565 => x"00000000",
   566 => x"00000000",
   567 => x"00000000",
   568 => x"00000000",
   569 => x"00000000",
   570 => x"00000000",
   571 => x"00000000",
   572 => x"00000888",
   573 => x"00000000",
   574 => x"00000000",
   575 => x"00000000",
   576 => x"00000000",
   577 => x"00000000",
   578 => x"00000000",
   579 => x"00000000",
   580 => x"00000000",
   581 => x"00000000",
   582 => x"00000000",
   583 => x"00000000",
   584 => x"00000000",
   585 => x"00000000",
   586 => x"00000000",
   587 => x"00000000",
   588 => x"00000000",
   589 => x"00000000",
   590 => x"00000000",
   591 => x"00000000",
   592 => x"00000000",
   593 => x"00000000",
   594 => x"00000000",
   595 => x"00000000",
   596 => x"00000000",
   597 => x"00000000",
   598 => x"00000000",
   599 => x"00000000",
   600 => x"00000000",
   601 => x"00000001",
   602 => x"330eabcd",
   603 => x"1234e66d",
   604 => x"deec0005",
   605 => x"000b0000",
   606 => x"00000000",
   607 => x"00000000",
   608 => x"00000000",
   609 => x"00000000",
   610 => x"00000000",
   611 => x"00000000",
   612 => x"00000000",
   613 => x"00000000",
   614 => x"00000000",
   615 => x"00000000",
   616 => x"00000000",
   617 => x"00000000",
   618 => x"00000000",
   619 => x"00000000",
   620 => x"00000000",
   621 => x"00000000",
   622 => x"00000000",
   623 => x"00000000",
   624 => x"00000000",
   625 => x"00000000",
   626 => x"00000000",
   627 => x"00000000",
   628 => x"00000000",
   629 => x"00000000",
   630 => x"00000000",
   631 => x"00000000",
   632 => x"00000000",
   633 => x"00000000",
   634 => x"00000000",
   635 => x"00000000",
   636 => x"00000000",
   637 => x"00000000",
   638 => x"00000000",
   639 => x"00000000",
   640 => x"00000000",
   641 => x"00000000",
   642 => x"00000000",
   643 => x"00000000",
   644 => x"00000000",
   645 => x"00000000",
   646 => x"00000000",
   647 => x"00000000",
   648 => x"00000000",
   649 => x"00000000",
   650 => x"00000000",
   651 => x"00000000",
   652 => x"00000000",
   653 => x"00000000",
   654 => x"00000000",
   655 => x"00000000",
   656 => x"00000000",
   657 => x"00000000",
   658 => x"00000000",
   659 => x"00000000",
   660 => x"00000000",
   661 => x"00000000",
   662 => x"00000000",
   663 => x"00000000",
   664 => x"00000000",
   665 => x"00000000",
   666 => x"00000000",
   667 => x"00000000",
   668 => x"00000000",
   669 => x"00000000",
   670 => x"00000000",
   671 => x"00000000",
   672 => x"00000000",
   673 => x"00000000",
   674 => x"00000000",
   675 => x"00000000",
   676 => x"00000000",
   677 => x"00000000",
   678 => x"00000000",
   679 => x"00000000",
   680 => x"00000000",
   681 => x"00000000",
   682 => x"00000000",
   683 => x"00000000",
   684 => x"00000000",
   685 => x"00000000",
   686 => x"00000000",
   687 => x"00000000",
   688 => x"00000000",
   689 => x"00000000",
   690 => x"00000000",
   691 => x"00000000",
   692 => x"00000000",
   693 => x"00000000",
   694 => x"00000000",
   695 => x"00000000",
   696 => x"00000000",
   697 => x"00000000",
   698 => x"00000000",
   699 => x"00000000",
   700 => x"00000000",
   701 => x"00000000",
   702 => x"00000000",
   703 => x"00000000",
   704 => x"00000000",
   705 => x"00000000",
   706 => x"00000000",
   707 => x"00000000",
   708 => x"00000000",
   709 => x"00000000",
   710 => x"00000000",
   711 => x"00000000",
   712 => x"00000000",
   713 => x"00000000",
   714 => x"00000000",
   715 => x"00000000",
   716 => x"00000000",
   717 => x"00000000",
   718 => x"00000000",
   719 => x"00000000",
   720 => x"00000000",
   721 => x"00000000",
   722 => x"00000000",
   723 => x"00000000",
   724 => x"00000000",
   725 => x"00000000",
   726 => x"00000000",
   727 => x"00000000",
   728 => x"00000000",
   729 => x"00000000",
   730 => x"00000000",
   731 => x"00000000",
   732 => x"00000000",
   733 => x"00000000",
   734 => x"00000000",
   735 => x"00000000",
   736 => x"00000000",
   737 => x"00000000",
   738 => x"00000000",
   739 => x"00000000",
   740 => x"00000000",
   741 => x"00000000",
   742 => x"00000000",
   743 => x"00000000",
   744 => x"00000000",
   745 => x"00000000",
   746 => x"00000000",
   747 => x"00000000",
   748 => x"00000000",
   749 => x"00000000",
   750 => x"00000000",
   751 => x"00000000",
   752 => x"00000000",
   753 => x"00000000",
   754 => x"00000000",
   755 => x"00000000",
   756 => x"00000000",
   757 => x"00000000",
   758 => x"00000000",
   759 => x"00000000",
   760 => x"00000000",
   761 => x"00000000",
   762 => x"00000000",
   763 => x"00000000",
   764 => x"00000000",
   765 => x"00000000",
   766 => x"00000000",
   767 => x"00000000",
   768 => x"00000000",
   769 => x"00000000",
   770 => x"00000000",
   771 => x"00000000",
   772 => x"00000000",
   773 => x"00000000",
   774 => x"00000000",
   775 => x"00000000",
   776 => x"00000000",
   777 => x"00000000",
   778 => x"00000000",
   779 => x"00000000",
   780 => x"00000000",
   781 => x"00000000",
   782 => x"ffffffff",
   783 => x"00000000",
   784 => x"ffffffff",
   785 => x"00000000",
   786 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
